magic
tech sky130A
magscale 1 2
timestamp 1654782658
<< obsli1 >>
rect 1104 2159 63664 64753
<< obsm1 >>
rect 14 1436 64754 64784
<< metal2 >>
rect 294 66185 350 66985
rect 846 66185 902 66985
rect 1398 66185 1454 66985
rect 1950 66185 2006 66985
rect 2502 66185 2558 66985
rect 3054 66185 3110 66985
rect 3698 66185 3754 66985
rect 4250 66185 4306 66985
rect 4802 66185 4858 66985
rect 5354 66185 5410 66985
rect 5906 66185 5962 66985
rect 6550 66185 6606 66985
rect 7102 66185 7158 66985
rect 7654 66185 7710 66985
rect 8206 66185 8262 66985
rect 8758 66185 8814 66985
rect 9310 66185 9366 66985
rect 9954 66185 10010 66985
rect 10506 66185 10562 66985
rect 11058 66185 11114 66985
rect 11610 66185 11666 66985
rect 12162 66185 12218 66985
rect 12806 66185 12862 66985
rect 13358 66185 13414 66985
rect 13910 66185 13966 66985
rect 14462 66185 14518 66985
rect 15014 66185 15070 66985
rect 15566 66185 15622 66985
rect 16210 66185 16266 66985
rect 16762 66185 16818 66985
rect 17314 66185 17370 66985
rect 17866 66185 17922 66985
rect 18418 66185 18474 66985
rect 19062 66185 19118 66985
rect 19614 66185 19670 66985
rect 20166 66185 20222 66985
rect 20718 66185 20774 66985
rect 21270 66185 21326 66985
rect 21914 66185 21970 66985
rect 22466 66185 22522 66985
rect 23018 66185 23074 66985
rect 23570 66185 23626 66985
rect 24122 66185 24178 66985
rect 24674 66185 24730 66985
rect 25318 66185 25374 66985
rect 25870 66185 25926 66985
rect 26422 66185 26478 66985
rect 26974 66185 27030 66985
rect 27526 66185 27582 66985
rect 28170 66185 28226 66985
rect 28722 66185 28778 66985
rect 29274 66185 29330 66985
rect 29826 66185 29882 66985
rect 30378 66185 30434 66985
rect 30930 66185 30986 66985
rect 31574 66185 31630 66985
rect 32126 66185 32182 66985
rect 32678 66185 32734 66985
rect 33230 66185 33286 66985
rect 33782 66185 33838 66985
rect 34426 66185 34482 66985
rect 34978 66185 35034 66985
rect 35530 66185 35586 66985
rect 36082 66185 36138 66985
rect 36634 66185 36690 66985
rect 37186 66185 37242 66985
rect 37830 66185 37886 66985
rect 38382 66185 38438 66985
rect 38934 66185 38990 66985
rect 39486 66185 39542 66985
rect 40038 66185 40094 66985
rect 40682 66185 40738 66985
rect 41234 66185 41290 66985
rect 41786 66185 41842 66985
rect 42338 66185 42394 66985
rect 42890 66185 42946 66985
rect 43534 66185 43590 66985
rect 44086 66185 44142 66985
rect 44638 66185 44694 66985
rect 45190 66185 45246 66985
rect 45742 66185 45798 66985
rect 46294 66185 46350 66985
rect 46938 66185 46994 66985
rect 47490 66185 47546 66985
rect 48042 66185 48098 66985
rect 48594 66185 48650 66985
rect 49146 66185 49202 66985
rect 49790 66185 49846 66985
rect 50342 66185 50398 66985
rect 50894 66185 50950 66985
rect 51446 66185 51502 66985
rect 51998 66185 52054 66985
rect 52550 66185 52606 66985
rect 53194 66185 53250 66985
rect 53746 66185 53802 66985
rect 54298 66185 54354 66985
rect 54850 66185 54906 66985
rect 55402 66185 55458 66985
rect 56046 66185 56102 66985
rect 56598 66185 56654 66985
rect 57150 66185 57206 66985
rect 57702 66185 57758 66985
rect 58254 66185 58310 66985
rect 58806 66185 58862 66985
rect 59450 66185 59506 66985
rect 60002 66185 60058 66985
rect 60554 66185 60610 66985
rect 61106 66185 61162 66985
rect 61658 66185 61714 66985
rect 62302 66185 62358 66985
rect 62854 66185 62910 66985
rect 63406 66185 63462 66985
rect 63958 66185 64014 66985
rect 64510 66185 64566 66985
rect 18 0 74 800
rect 110 0 166 800
rect 202 0 258 800
rect 386 0 442 800
rect 478 0 534 800
rect 662 0 718 800
rect 754 0 810 800
rect 938 0 994 800
rect 1030 0 1086 800
rect 1122 0 1178 800
rect 1306 0 1362 800
rect 1398 0 1454 800
rect 1582 0 1638 800
rect 1674 0 1730 800
rect 1858 0 1914 800
rect 1950 0 2006 800
rect 2042 0 2098 800
rect 2226 0 2282 800
rect 2318 0 2374 800
rect 2502 0 2558 800
rect 2594 0 2650 800
rect 2778 0 2834 800
rect 2870 0 2926 800
rect 2962 0 3018 800
rect 3146 0 3202 800
rect 3238 0 3294 800
rect 3422 0 3478 800
rect 3514 0 3570 800
rect 3698 0 3754 800
rect 3790 0 3846 800
rect 3882 0 3938 800
rect 4066 0 4122 800
rect 4158 0 4214 800
rect 4342 0 4398 800
rect 4434 0 4490 800
rect 4618 0 4674 800
rect 4710 0 4766 800
rect 4802 0 4858 800
rect 4986 0 5042 800
rect 5078 0 5134 800
rect 5262 0 5318 800
rect 5354 0 5410 800
rect 5538 0 5594 800
rect 5630 0 5686 800
rect 5722 0 5778 800
rect 5906 0 5962 800
rect 5998 0 6054 800
rect 6182 0 6238 800
rect 6274 0 6330 800
rect 6458 0 6514 800
rect 6550 0 6606 800
rect 6642 0 6698 800
rect 6826 0 6882 800
rect 6918 0 6974 800
rect 7102 0 7158 800
rect 7194 0 7250 800
rect 7378 0 7434 800
rect 7470 0 7526 800
rect 7562 0 7618 800
rect 7746 0 7802 800
rect 7838 0 7894 800
rect 8022 0 8078 800
rect 8114 0 8170 800
rect 8298 0 8354 800
rect 8390 0 8446 800
rect 8482 0 8538 800
rect 8666 0 8722 800
rect 8758 0 8814 800
rect 8942 0 8998 800
rect 9034 0 9090 800
rect 9218 0 9274 800
rect 9310 0 9366 800
rect 9402 0 9458 800
rect 9586 0 9642 800
rect 9678 0 9734 800
rect 9862 0 9918 800
rect 9954 0 10010 800
rect 10138 0 10194 800
rect 10230 0 10286 800
rect 10322 0 10378 800
rect 10506 0 10562 800
rect 10598 0 10654 800
rect 10782 0 10838 800
rect 10874 0 10930 800
rect 11058 0 11114 800
rect 11150 0 11206 800
rect 11242 0 11298 800
rect 11426 0 11482 800
rect 11518 0 11574 800
rect 11702 0 11758 800
rect 11794 0 11850 800
rect 11978 0 12034 800
rect 12070 0 12126 800
rect 12162 0 12218 800
rect 12346 0 12402 800
rect 12438 0 12494 800
rect 12622 0 12678 800
rect 12714 0 12770 800
rect 12898 0 12954 800
rect 12990 0 13046 800
rect 13174 0 13230 800
rect 13266 0 13322 800
rect 13358 0 13414 800
rect 13542 0 13598 800
rect 13634 0 13690 800
rect 13818 0 13874 800
rect 13910 0 13966 800
rect 14094 0 14150 800
rect 14186 0 14242 800
rect 14278 0 14334 800
rect 14462 0 14518 800
rect 14554 0 14610 800
rect 14738 0 14794 800
rect 14830 0 14886 800
rect 15014 0 15070 800
rect 15106 0 15162 800
rect 15198 0 15254 800
rect 15382 0 15438 800
rect 15474 0 15530 800
rect 15658 0 15714 800
rect 15750 0 15806 800
rect 15934 0 15990 800
rect 16026 0 16082 800
rect 16118 0 16174 800
rect 16302 0 16358 800
rect 16394 0 16450 800
rect 16578 0 16634 800
rect 16670 0 16726 800
rect 16854 0 16910 800
rect 16946 0 17002 800
rect 17038 0 17094 800
rect 17222 0 17278 800
rect 17314 0 17370 800
rect 17498 0 17554 800
rect 17590 0 17646 800
rect 17774 0 17830 800
rect 17866 0 17922 800
rect 17958 0 18014 800
rect 18142 0 18198 800
rect 18234 0 18290 800
rect 18418 0 18474 800
rect 18510 0 18566 800
rect 18694 0 18750 800
rect 18786 0 18842 800
rect 18878 0 18934 800
rect 19062 0 19118 800
rect 19154 0 19210 800
rect 19338 0 19394 800
rect 19430 0 19486 800
rect 19614 0 19670 800
rect 19706 0 19762 800
rect 19798 0 19854 800
rect 19982 0 20038 800
rect 20074 0 20130 800
rect 20258 0 20314 800
rect 20350 0 20406 800
rect 20534 0 20590 800
rect 20626 0 20682 800
rect 20718 0 20774 800
rect 20902 0 20958 800
rect 20994 0 21050 800
rect 21178 0 21234 800
rect 21270 0 21326 800
rect 21454 0 21510 800
rect 21546 0 21602 800
rect 21638 0 21694 800
rect 21822 0 21878 800
rect 21914 0 21970 800
rect 22098 0 22154 800
rect 22190 0 22246 800
rect 22374 0 22430 800
rect 22466 0 22522 800
rect 22558 0 22614 800
rect 22742 0 22798 800
rect 22834 0 22890 800
rect 23018 0 23074 800
rect 23110 0 23166 800
rect 23294 0 23350 800
rect 23386 0 23442 800
rect 23478 0 23534 800
rect 23662 0 23718 800
rect 23754 0 23810 800
rect 23938 0 23994 800
rect 24030 0 24086 800
rect 24214 0 24270 800
rect 24306 0 24362 800
rect 24398 0 24454 800
rect 24582 0 24638 800
rect 24674 0 24730 800
rect 24858 0 24914 800
rect 24950 0 25006 800
rect 25134 0 25190 800
rect 25226 0 25282 800
rect 25318 0 25374 800
rect 25502 0 25558 800
rect 25594 0 25650 800
rect 25778 0 25834 800
rect 25870 0 25926 800
rect 26054 0 26110 800
rect 26146 0 26202 800
rect 26330 0 26386 800
rect 26422 0 26478 800
rect 26514 0 26570 800
rect 26698 0 26754 800
rect 26790 0 26846 800
rect 26974 0 27030 800
rect 27066 0 27122 800
rect 27250 0 27306 800
rect 27342 0 27398 800
rect 27434 0 27490 800
rect 27618 0 27674 800
rect 27710 0 27766 800
rect 27894 0 27950 800
rect 27986 0 28042 800
rect 28170 0 28226 800
rect 28262 0 28318 800
rect 28354 0 28410 800
rect 28538 0 28594 800
rect 28630 0 28686 800
rect 28814 0 28870 800
rect 28906 0 28962 800
rect 29090 0 29146 800
rect 29182 0 29238 800
rect 29274 0 29330 800
rect 29458 0 29514 800
rect 29550 0 29606 800
rect 29734 0 29790 800
rect 29826 0 29882 800
rect 30010 0 30066 800
rect 30102 0 30158 800
rect 30194 0 30250 800
rect 30378 0 30434 800
rect 30470 0 30526 800
rect 30654 0 30710 800
rect 30746 0 30802 800
rect 30930 0 30986 800
rect 31022 0 31078 800
rect 31114 0 31170 800
rect 31298 0 31354 800
rect 31390 0 31446 800
rect 31574 0 31630 800
rect 31666 0 31722 800
rect 31850 0 31906 800
rect 31942 0 31998 800
rect 32034 0 32090 800
rect 32218 0 32274 800
rect 32310 0 32366 800
rect 32494 0 32550 800
rect 32586 0 32642 800
rect 32770 0 32826 800
rect 32862 0 32918 800
rect 32954 0 33010 800
rect 33138 0 33194 800
rect 33230 0 33286 800
rect 33414 0 33470 800
rect 33506 0 33562 800
rect 33690 0 33746 800
rect 33782 0 33838 800
rect 33874 0 33930 800
rect 34058 0 34114 800
rect 34150 0 34206 800
rect 34334 0 34390 800
rect 34426 0 34482 800
rect 34610 0 34666 800
rect 34702 0 34758 800
rect 34794 0 34850 800
rect 34978 0 35034 800
rect 35070 0 35126 800
rect 35254 0 35310 800
rect 35346 0 35402 800
rect 35530 0 35586 800
rect 35622 0 35678 800
rect 35714 0 35770 800
rect 35898 0 35954 800
rect 35990 0 36046 800
rect 36174 0 36230 800
rect 36266 0 36322 800
rect 36450 0 36506 800
rect 36542 0 36598 800
rect 36634 0 36690 800
rect 36818 0 36874 800
rect 36910 0 36966 800
rect 37094 0 37150 800
rect 37186 0 37242 800
rect 37370 0 37426 800
rect 37462 0 37518 800
rect 37554 0 37610 800
rect 37738 0 37794 800
rect 37830 0 37886 800
rect 38014 0 38070 800
rect 38106 0 38162 800
rect 38290 0 38346 800
rect 38382 0 38438 800
rect 38474 0 38530 800
rect 38658 0 38714 800
rect 38750 0 38806 800
rect 38934 0 38990 800
rect 39026 0 39082 800
rect 39210 0 39266 800
rect 39302 0 39358 800
rect 39486 0 39542 800
rect 39578 0 39634 800
rect 39670 0 39726 800
rect 39854 0 39910 800
rect 39946 0 40002 800
rect 40130 0 40186 800
rect 40222 0 40278 800
rect 40406 0 40462 800
rect 40498 0 40554 800
rect 40590 0 40646 800
rect 40774 0 40830 800
rect 40866 0 40922 800
rect 41050 0 41106 800
rect 41142 0 41198 800
rect 41326 0 41382 800
rect 41418 0 41474 800
rect 41510 0 41566 800
rect 41694 0 41750 800
rect 41786 0 41842 800
rect 41970 0 42026 800
rect 42062 0 42118 800
rect 42246 0 42302 800
rect 42338 0 42394 800
rect 42430 0 42486 800
rect 42614 0 42670 800
rect 42706 0 42762 800
rect 42890 0 42946 800
rect 42982 0 43038 800
rect 43166 0 43222 800
rect 43258 0 43314 800
rect 43350 0 43406 800
rect 43534 0 43590 800
rect 43626 0 43682 800
rect 43810 0 43866 800
rect 43902 0 43958 800
rect 44086 0 44142 800
rect 44178 0 44234 800
rect 44270 0 44326 800
rect 44454 0 44510 800
rect 44546 0 44602 800
rect 44730 0 44786 800
rect 44822 0 44878 800
rect 45006 0 45062 800
rect 45098 0 45154 800
rect 45190 0 45246 800
rect 45374 0 45430 800
rect 45466 0 45522 800
rect 45650 0 45706 800
rect 45742 0 45798 800
rect 45926 0 45982 800
rect 46018 0 46074 800
rect 46110 0 46166 800
rect 46294 0 46350 800
rect 46386 0 46442 800
rect 46570 0 46626 800
rect 46662 0 46718 800
rect 46846 0 46902 800
rect 46938 0 46994 800
rect 47030 0 47086 800
rect 47214 0 47270 800
rect 47306 0 47362 800
rect 47490 0 47546 800
rect 47582 0 47638 800
rect 47766 0 47822 800
rect 47858 0 47914 800
rect 47950 0 48006 800
rect 48134 0 48190 800
rect 48226 0 48282 800
rect 48410 0 48466 800
rect 48502 0 48558 800
rect 48686 0 48742 800
rect 48778 0 48834 800
rect 48870 0 48926 800
rect 49054 0 49110 800
rect 49146 0 49202 800
rect 49330 0 49386 800
rect 49422 0 49478 800
rect 49606 0 49662 800
rect 49698 0 49754 800
rect 49790 0 49846 800
rect 49974 0 50030 800
rect 50066 0 50122 800
rect 50250 0 50306 800
rect 50342 0 50398 800
rect 50526 0 50582 800
rect 50618 0 50674 800
rect 50710 0 50766 800
rect 50894 0 50950 800
rect 50986 0 51042 800
rect 51170 0 51226 800
rect 51262 0 51318 800
rect 51446 0 51502 800
rect 51538 0 51594 800
rect 51630 0 51686 800
rect 51814 0 51870 800
rect 51906 0 51962 800
rect 52090 0 52146 800
rect 52182 0 52238 800
rect 52366 0 52422 800
rect 52458 0 52514 800
rect 52642 0 52698 800
rect 52734 0 52790 800
rect 52826 0 52882 800
rect 53010 0 53066 800
rect 53102 0 53158 800
rect 53286 0 53342 800
rect 53378 0 53434 800
rect 53562 0 53618 800
rect 53654 0 53710 800
rect 53746 0 53802 800
rect 53930 0 53986 800
rect 54022 0 54078 800
rect 54206 0 54262 800
rect 54298 0 54354 800
rect 54482 0 54538 800
rect 54574 0 54630 800
rect 54666 0 54722 800
rect 54850 0 54906 800
rect 54942 0 54998 800
rect 55126 0 55182 800
rect 55218 0 55274 800
rect 55402 0 55458 800
rect 55494 0 55550 800
rect 55586 0 55642 800
rect 55770 0 55826 800
rect 55862 0 55918 800
rect 56046 0 56102 800
rect 56138 0 56194 800
rect 56322 0 56378 800
rect 56414 0 56470 800
rect 56506 0 56562 800
rect 56690 0 56746 800
rect 56782 0 56838 800
rect 56966 0 57022 800
rect 57058 0 57114 800
rect 57242 0 57298 800
rect 57334 0 57390 800
rect 57426 0 57482 800
rect 57610 0 57666 800
rect 57702 0 57758 800
rect 57886 0 57942 800
rect 57978 0 58034 800
rect 58162 0 58218 800
rect 58254 0 58310 800
rect 58346 0 58402 800
rect 58530 0 58586 800
rect 58622 0 58678 800
rect 58806 0 58862 800
rect 58898 0 58954 800
rect 59082 0 59138 800
rect 59174 0 59230 800
rect 59266 0 59322 800
rect 59450 0 59506 800
rect 59542 0 59598 800
rect 59726 0 59782 800
rect 59818 0 59874 800
rect 60002 0 60058 800
rect 60094 0 60150 800
rect 60186 0 60242 800
rect 60370 0 60426 800
rect 60462 0 60518 800
rect 60646 0 60702 800
rect 60738 0 60794 800
rect 60922 0 60978 800
rect 61014 0 61070 800
rect 61106 0 61162 800
rect 61290 0 61346 800
rect 61382 0 61438 800
rect 61566 0 61622 800
rect 61658 0 61714 800
rect 61842 0 61898 800
rect 61934 0 61990 800
rect 62026 0 62082 800
rect 62210 0 62266 800
rect 62302 0 62358 800
rect 62486 0 62542 800
rect 62578 0 62634 800
rect 62762 0 62818 800
rect 62854 0 62910 800
rect 62946 0 63002 800
rect 63130 0 63186 800
rect 63222 0 63278 800
rect 63406 0 63462 800
rect 63498 0 63554 800
rect 63682 0 63738 800
rect 63774 0 63830 800
rect 63866 0 63922 800
rect 64050 0 64106 800
rect 64142 0 64198 800
rect 64326 0 64382 800
rect 64418 0 64474 800
rect 64602 0 64658 800
rect 64694 0 64750 800
<< obsm2 >>
rect 20 66129 238 66314
rect 406 66129 790 66314
rect 958 66129 1342 66314
rect 1510 66129 1894 66314
rect 2062 66129 2446 66314
rect 2614 66129 2998 66314
rect 3166 66129 3642 66314
rect 3810 66129 4194 66314
rect 4362 66129 4746 66314
rect 4914 66129 5298 66314
rect 5466 66129 5850 66314
rect 6018 66129 6494 66314
rect 6662 66129 7046 66314
rect 7214 66129 7598 66314
rect 7766 66129 8150 66314
rect 8318 66129 8702 66314
rect 8870 66129 9254 66314
rect 9422 66129 9898 66314
rect 10066 66129 10450 66314
rect 10618 66129 11002 66314
rect 11170 66129 11554 66314
rect 11722 66129 12106 66314
rect 12274 66129 12750 66314
rect 12918 66129 13302 66314
rect 13470 66129 13854 66314
rect 14022 66129 14406 66314
rect 14574 66129 14958 66314
rect 15126 66129 15510 66314
rect 15678 66129 16154 66314
rect 16322 66129 16706 66314
rect 16874 66129 17258 66314
rect 17426 66129 17810 66314
rect 17978 66129 18362 66314
rect 18530 66129 19006 66314
rect 19174 66129 19558 66314
rect 19726 66129 20110 66314
rect 20278 66129 20662 66314
rect 20830 66129 21214 66314
rect 21382 66129 21858 66314
rect 22026 66129 22410 66314
rect 22578 66129 22962 66314
rect 23130 66129 23514 66314
rect 23682 66129 24066 66314
rect 24234 66129 24618 66314
rect 24786 66129 25262 66314
rect 25430 66129 25814 66314
rect 25982 66129 26366 66314
rect 26534 66129 26918 66314
rect 27086 66129 27470 66314
rect 27638 66129 28114 66314
rect 28282 66129 28666 66314
rect 28834 66129 29218 66314
rect 29386 66129 29770 66314
rect 29938 66129 30322 66314
rect 30490 66129 30874 66314
rect 31042 66129 31518 66314
rect 31686 66129 32070 66314
rect 32238 66129 32622 66314
rect 32790 66129 33174 66314
rect 33342 66129 33726 66314
rect 33894 66129 34370 66314
rect 34538 66129 34922 66314
rect 35090 66129 35474 66314
rect 35642 66129 36026 66314
rect 36194 66129 36578 66314
rect 36746 66129 37130 66314
rect 37298 66129 37774 66314
rect 37942 66129 38326 66314
rect 38494 66129 38878 66314
rect 39046 66129 39430 66314
rect 39598 66129 39982 66314
rect 40150 66129 40626 66314
rect 40794 66129 41178 66314
rect 41346 66129 41730 66314
rect 41898 66129 42282 66314
rect 42450 66129 42834 66314
rect 43002 66129 43478 66314
rect 43646 66129 44030 66314
rect 44198 66129 44582 66314
rect 44750 66129 45134 66314
rect 45302 66129 45686 66314
rect 45854 66129 46238 66314
rect 46406 66129 46882 66314
rect 47050 66129 47434 66314
rect 47602 66129 47986 66314
rect 48154 66129 48538 66314
rect 48706 66129 49090 66314
rect 49258 66129 49734 66314
rect 49902 66129 50286 66314
rect 50454 66129 50838 66314
rect 51006 66129 51390 66314
rect 51558 66129 51942 66314
rect 52110 66129 52494 66314
rect 52662 66129 53138 66314
rect 53306 66129 53690 66314
rect 53858 66129 54242 66314
rect 54410 66129 54794 66314
rect 54962 66129 55346 66314
rect 55514 66129 55990 66314
rect 56158 66129 56542 66314
rect 56710 66129 57094 66314
rect 57262 66129 57646 66314
rect 57814 66129 58198 66314
rect 58366 66129 58750 66314
rect 58918 66129 59394 66314
rect 59562 66129 59946 66314
rect 60114 66129 60498 66314
rect 60666 66129 61050 66314
rect 61218 66129 61602 66314
rect 61770 66129 62246 66314
rect 62414 66129 62798 66314
rect 62966 66129 63350 66314
rect 63518 66129 63902 66314
rect 64070 66129 64454 66314
rect 64622 66129 64748 66314
rect 20 856 64748 66129
rect 314 800 330 856
rect 590 800 606 856
rect 866 800 882 856
rect 1234 800 1250 856
rect 1510 800 1526 856
rect 1786 800 1802 856
rect 2154 800 2170 856
rect 2430 800 2446 856
rect 2706 800 2722 856
rect 3074 800 3090 856
rect 3350 800 3366 856
rect 3626 800 3642 856
rect 3994 800 4010 856
rect 4270 800 4286 856
rect 4546 800 4562 856
rect 4914 800 4930 856
rect 5190 800 5206 856
rect 5466 800 5482 856
rect 5834 800 5850 856
rect 6110 800 6126 856
rect 6386 800 6402 856
rect 6754 800 6770 856
rect 7030 800 7046 856
rect 7306 800 7322 856
rect 7674 800 7690 856
rect 7950 800 7966 856
rect 8226 800 8242 856
rect 8594 800 8610 856
rect 8870 800 8886 856
rect 9146 800 9162 856
rect 9514 800 9530 856
rect 9790 800 9806 856
rect 10066 800 10082 856
rect 10434 800 10450 856
rect 10710 800 10726 856
rect 10986 800 11002 856
rect 11354 800 11370 856
rect 11630 800 11646 856
rect 11906 800 11922 856
rect 12274 800 12290 856
rect 12550 800 12566 856
rect 12826 800 12842 856
rect 13102 800 13118 856
rect 13470 800 13486 856
rect 13746 800 13762 856
rect 14022 800 14038 856
rect 14390 800 14406 856
rect 14666 800 14682 856
rect 14942 800 14958 856
rect 15310 800 15326 856
rect 15586 800 15602 856
rect 15862 800 15878 856
rect 16230 800 16246 856
rect 16506 800 16522 856
rect 16782 800 16798 856
rect 17150 800 17166 856
rect 17426 800 17442 856
rect 17702 800 17718 856
rect 18070 800 18086 856
rect 18346 800 18362 856
rect 18622 800 18638 856
rect 18990 800 19006 856
rect 19266 800 19282 856
rect 19542 800 19558 856
rect 19910 800 19926 856
rect 20186 800 20202 856
rect 20462 800 20478 856
rect 20830 800 20846 856
rect 21106 800 21122 856
rect 21382 800 21398 856
rect 21750 800 21766 856
rect 22026 800 22042 856
rect 22302 800 22318 856
rect 22670 800 22686 856
rect 22946 800 22962 856
rect 23222 800 23238 856
rect 23590 800 23606 856
rect 23866 800 23882 856
rect 24142 800 24158 856
rect 24510 800 24526 856
rect 24786 800 24802 856
rect 25062 800 25078 856
rect 25430 800 25446 856
rect 25706 800 25722 856
rect 25982 800 25998 856
rect 26258 800 26274 856
rect 26626 800 26642 856
rect 26902 800 26918 856
rect 27178 800 27194 856
rect 27546 800 27562 856
rect 27822 800 27838 856
rect 28098 800 28114 856
rect 28466 800 28482 856
rect 28742 800 28758 856
rect 29018 800 29034 856
rect 29386 800 29402 856
rect 29662 800 29678 856
rect 29938 800 29954 856
rect 30306 800 30322 856
rect 30582 800 30598 856
rect 30858 800 30874 856
rect 31226 800 31242 856
rect 31502 800 31518 856
rect 31778 800 31794 856
rect 32146 800 32162 856
rect 32422 800 32438 856
rect 32698 800 32714 856
rect 33066 800 33082 856
rect 33342 800 33358 856
rect 33618 800 33634 856
rect 33986 800 34002 856
rect 34262 800 34278 856
rect 34538 800 34554 856
rect 34906 800 34922 856
rect 35182 800 35198 856
rect 35458 800 35474 856
rect 35826 800 35842 856
rect 36102 800 36118 856
rect 36378 800 36394 856
rect 36746 800 36762 856
rect 37022 800 37038 856
rect 37298 800 37314 856
rect 37666 800 37682 856
rect 37942 800 37958 856
rect 38218 800 38234 856
rect 38586 800 38602 856
rect 38862 800 38878 856
rect 39138 800 39154 856
rect 39414 800 39430 856
rect 39782 800 39798 856
rect 40058 800 40074 856
rect 40334 800 40350 856
rect 40702 800 40718 856
rect 40978 800 40994 856
rect 41254 800 41270 856
rect 41622 800 41638 856
rect 41898 800 41914 856
rect 42174 800 42190 856
rect 42542 800 42558 856
rect 42818 800 42834 856
rect 43094 800 43110 856
rect 43462 800 43478 856
rect 43738 800 43754 856
rect 44014 800 44030 856
rect 44382 800 44398 856
rect 44658 800 44674 856
rect 44934 800 44950 856
rect 45302 800 45318 856
rect 45578 800 45594 856
rect 45854 800 45870 856
rect 46222 800 46238 856
rect 46498 800 46514 856
rect 46774 800 46790 856
rect 47142 800 47158 856
rect 47418 800 47434 856
rect 47694 800 47710 856
rect 48062 800 48078 856
rect 48338 800 48354 856
rect 48614 800 48630 856
rect 48982 800 48998 856
rect 49258 800 49274 856
rect 49534 800 49550 856
rect 49902 800 49918 856
rect 50178 800 50194 856
rect 50454 800 50470 856
rect 50822 800 50838 856
rect 51098 800 51114 856
rect 51374 800 51390 856
rect 51742 800 51758 856
rect 52018 800 52034 856
rect 52294 800 52310 856
rect 52570 800 52586 856
rect 52938 800 52954 856
rect 53214 800 53230 856
rect 53490 800 53506 856
rect 53858 800 53874 856
rect 54134 800 54150 856
rect 54410 800 54426 856
rect 54778 800 54794 856
rect 55054 800 55070 856
rect 55330 800 55346 856
rect 55698 800 55714 856
rect 55974 800 55990 856
rect 56250 800 56266 856
rect 56618 800 56634 856
rect 56894 800 56910 856
rect 57170 800 57186 856
rect 57538 800 57554 856
rect 57814 800 57830 856
rect 58090 800 58106 856
rect 58458 800 58474 856
rect 58734 800 58750 856
rect 59010 800 59026 856
rect 59378 800 59394 856
rect 59654 800 59670 856
rect 59930 800 59946 856
rect 60298 800 60314 856
rect 60574 800 60590 856
rect 60850 800 60866 856
rect 61218 800 61234 856
rect 61494 800 61510 856
rect 61770 800 61786 856
rect 62138 800 62154 856
rect 62414 800 62430 856
rect 62690 800 62706 856
rect 63058 800 63074 856
rect 63334 800 63350 856
rect 63610 800 63626 856
rect 63978 800 63994 856
rect 64254 800 64270 856
rect 64530 800 64546 856
<< obsm3 >>
rect 4208 2143 60799 64769
<< metal4 >>
rect 4208 2128 4528 64784
rect 19568 2128 19888 64784
rect 34928 2128 35248 64784
rect 50288 2128 50608 64784
<< obsm4 >>
rect 20851 11867 34848 64429
rect 35328 11867 47229 64429
<< labels >>
rlabel metal2 s 294 66185 350 66985 6 io_in[0]
port 1 nsew signal input
rlabel metal2 s 17314 66185 17370 66985 6 io_in[10]
port 2 nsew signal input
rlabel metal2 s 19062 66185 19118 66985 6 io_in[11]
port 3 nsew signal input
rlabel metal2 s 20718 66185 20774 66985 6 io_in[12]
port 4 nsew signal input
rlabel metal2 s 22466 66185 22522 66985 6 io_in[13]
port 5 nsew signal input
rlabel metal2 s 24122 66185 24178 66985 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 25870 66185 25926 66985 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 27526 66185 27582 66985 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 29274 66185 29330 66985 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 30930 66185 30986 66985 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 32678 66185 32734 66985 6 io_in[19]
port 11 nsew signal input
rlabel metal2 s 1950 66185 2006 66985 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 34426 66185 34482 66985 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 36082 66185 36138 66985 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 37830 66185 37886 66985 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 39486 66185 39542 66985 6 io_in[23]
port 16 nsew signal input
rlabel metal2 s 41234 66185 41290 66985 6 io_in[24]
port 17 nsew signal input
rlabel metal2 s 42890 66185 42946 66985 6 io_in[25]
port 18 nsew signal input
rlabel metal2 s 44638 66185 44694 66985 6 io_in[26]
port 19 nsew signal input
rlabel metal2 s 46294 66185 46350 66985 6 io_in[27]
port 20 nsew signal input
rlabel metal2 s 48042 66185 48098 66985 6 io_in[28]
port 21 nsew signal input
rlabel metal2 s 49790 66185 49846 66985 6 io_in[29]
port 22 nsew signal input
rlabel metal2 s 3698 66185 3754 66985 6 io_in[2]
port 23 nsew signal input
rlabel metal2 s 51446 66185 51502 66985 6 io_in[30]
port 24 nsew signal input
rlabel metal2 s 53194 66185 53250 66985 6 io_in[31]
port 25 nsew signal input
rlabel metal2 s 54850 66185 54906 66985 6 io_in[32]
port 26 nsew signal input
rlabel metal2 s 56598 66185 56654 66985 6 io_in[33]
port 27 nsew signal input
rlabel metal2 s 58254 66185 58310 66985 6 io_in[34]
port 28 nsew signal input
rlabel metal2 s 60002 66185 60058 66985 6 io_in[35]
port 29 nsew signal input
rlabel metal2 s 61658 66185 61714 66985 6 io_in[36]
port 30 nsew signal input
rlabel metal2 s 63406 66185 63462 66985 6 io_in[37]
port 31 nsew signal input
rlabel metal2 s 5354 66185 5410 66985 6 io_in[3]
port 32 nsew signal input
rlabel metal2 s 7102 66185 7158 66985 6 io_in[4]
port 33 nsew signal input
rlabel metal2 s 8758 66185 8814 66985 6 io_in[5]
port 34 nsew signal input
rlabel metal2 s 10506 66185 10562 66985 6 io_in[6]
port 35 nsew signal input
rlabel metal2 s 12162 66185 12218 66985 6 io_in[7]
port 36 nsew signal input
rlabel metal2 s 13910 66185 13966 66985 6 io_in[8]
port 37 nsew signal input
rlabel metal2 s 15566 66185 15622 66985 6 io_in[9]
port 38 nsew signal input
rlabel metal2 s 846 66185 902 66985 6 io_oeb[0]
port 39 nsew signal output
rlabel metal2 s 17866 66185 17922 66985 6 io_oeb[10]
port 40 nsew signal output
rlabel metal2 s 19614 66185 19670 66985 6 io_oeb[11]
port 41 nsew signal output
rlabel metal2 s 21270 66185 21326 66985 6 io_oeb[12]
port 42 nsew signal output
rlabel metal2 s 23018 66185 23074 66985 6 io_oeb[13]
port 43 nsew signal output
rlabel metal2 s 24674 66185 24730 66985 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 26422 66185 26478 66985 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 28170 66185 28226 66985 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 29826 66185 29882 66985 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 31574 66185 31630 66985 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 33230 66185 33286 66985 6 io_oeb[19]
port 49 nsew signal output
rlabel metal2 s 2502 66185 2558 66985 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 34978 66185 35034 66985 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 36634 66185 36690 66985 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 38382 66185 38438 66985 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 40038 66185 40094 66985 6 io_oeb[23]
port 54 nsew signal output
rlabel metal2 s 41786 66185 41842 66985 6 io_oeb[24]
port 55 nsew signal output
rlabel metal2 s 43534 66185 43590 66985 6 io_oeb[25]
port 56 nsew signal output
rlabel metal2 s 45190 66185 45246 66985 6 io_oeb[26]
port 57 nsew signal output
rlabel metal2 s 46938 66185 46994 66985 6 io_oeb[27]
port 58 nsew signal output
rlabel metal2 s 48594 66185 48650 66985 6 io_oeb[28]
port 59 nsew signal output
rlabel metal2 s 50342 66185 50398 66985 6 io_oeb[29]
port 60 nsew signal output
rlabel metal2 s 4250 66185 4306 66985 6 io_oeb[2]
port 61 nsew signal output
rlabel metal2 s 51998 66185 52054 66985 6 io_oeb[30]
port 62 nsew signal output
rlabel metal2 s 53746 66185 53802 66985 6 io_oeb[31]
port 63 nsew signal output
rlabel metal2 s 55402 66185 55458 66985 6 io_oeb[32]
port 64 nsew signal output
rlabel metal2 s 57150 66185 57206 66985 6 io_oeb[33]
port 65 nsew signal output
rlabel metal2 s 58806 66185 58862 66985 6 io_oeb[34]
port 66 nsew signal output
rlabel metal2 s 60554 66185 60610 66985 6 io_oeb[35]
port 67 nsew signal output
rlabel metal2 s 62302 66185 62358 66985 6 io_oeb[36]
port 68 nsew signal output
rlabel metal2 s 63958 66185 64014 66985 6 io_oeb[37]
port 69 nsew signal output
rlabel metal2 s 5906 66185 5962 66985 6 io_oeb[3]
port 70 nsew signal output
rlabel metal2 s 7654 66185 7710 66985 6 io_oeb[4]
port 71 nsew signal output
rlabel metal2 s 9310 66185 9366 66985 6 io_oeb[5]
port 72 nsew signal output
rlabel metal2 s 11058 66185 11114 66985 6 io_oeb[6]
port 73 nsew signal output
rlabel metal2 s 12806 66185 12862 66985 6 io_oeb[7]
port 74 nsew signal output
rlabel metal2 s 14462 66185 14518 66985 6 io_oeb[8]
port 75 nsew signal output
rlabel metal2 s 16210 66185 16266 66985 6 io_oeb[9]
port 76 nsew signal output
rlabel metal2 s 1398 66185 1454 66985 6 io_out[0]
port 77 nsew signal output
rlabel metal2 s 18418 66185 18474 66985 6 io_out[10]
port 78 nsew signal output
rlabel metal2 s 20166 66185 20222 66985 6 io_out[11]
port 79 nsew signal output
rlabel metal2 s 21914 66185 21970 66985 6 io_out[12]
port 80 nsew signal output
rlabel metal2 s 23570 66185 23626 66985 6 io_out[13]
port 81 nsew signal output
rlabel metal2 s 25318 66185 25374 66985 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 26974 66185 27030 66985 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 28722 66185 28778 66985 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 30378 66185 30434 66985 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 32126 66185 32182 66985 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 33782 66185 33838 66985 6 io_out[19]
port 87 nsew signal output
rlabel metal2 s 3054 66185 3110 66985 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 35530 66185 35586 66985 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 37186 66185 37242 66985 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 38934 66185 38990 66985 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 40682 66185 40738 66985 6 io_out[23]
port 92 nsew signal output
rlabel metal2 s 42338 66185 42394 66985 6 io_out[24]
port 93 nsew signal output
rlabel metal2 s 44086 66185 44142 66985 6 io_out[25]
port 94 nsew signal output
rlabel metal2 s 45742 66185 45798 66985 6 io_out[26]
port 95 nsew signal output
rlabel metal2 s 47490 66185 47546 66985 6 io_out[27]
port 96 nsew signal output
rlabel metal2 s 49146 66185 49202 66985 6 io_out[28]
port 97 nsew signal output
rlabel metal2 s 50894 66185 50950 66985 6 io_out[29]
port 98 nsew signal output
rlabel metal2 s 4802 66185 4858 66985 6 io_out[2]
port 99 nsew signal output
rlabel metal2 s 52550 66185 52606 66985 6 io_out[30]
port 100 nsew signal output
rlabel metal2 s 54298 66185 54354 66985 6 io_out[31]
port 101 nsew signal output
rlabel metal2 s 56046 66185 56102 66985 6 io_out[32]
port 102 nsew signal output
rlabel metal2 s 57702 66185 57758 66985 6 io_out[33]
port 103 nsew signal output
rlabel metal2 s 59450 66185 59506 66985 6 io_out[34]
port 104 nsew signal output
rlabel metal2 s 61106 66185 61162 66985 6 io_out[35]
port 105 nsew signal output
rlabel metal2 s 62854 66185 62910 66985 6 io_out[36]
port 106 nsew signal output
rlabel metal2 s 64510 66185 64566 66985 6 io_out[37]
port 107 nsew signal output
rlabel metal2 s 6550 66185 6606 66985 6 io_out[3]
port 108 nsew signal output
rlabel metal2 s 8206 66185 8262 66985 6 io_out[4]
port 109 nsew signal output
rlabel metal2 s 9954 66185 10010 66985 6 io_out[5]
port 110 nsew signal output
rlabel metal2 s 11610 66185 11666 66985 6 io_out[6]
port 111 nsew signal output
rlabel metal2 s 13358 66185 13414 66985 6 io_out[7]
port 112 nsew signal output
rlabel metal2 s 15014 66185 15070 66985 6 io_out[8]
port 113 nsew signal output
rlabel metal2 s 16762 66185 16818 66985 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 64418 0 64474 800 6 irq[0]
port 115 nsew signal output
rlabel metal2 s 64602 0 64658 800 6 irq[1]
port 116 nsew signal output
rlabel metal2 s 64694 0 64750 800 6 irq[2]
port 117 nsew signal output
rlabel metal2 s 13910 0 13966 800 6 la_data_in[0]
port 118 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[100]
port 119 nsew signal input
rlabel metal2 s 53746 0 53802 800 6 la_data_in[101]
port 120 nsew signal input
rlabel metal2 s 54206 0 54262 800 6 la_data_in[102]
port 121 nsew signal input
rlabel metal2 s 54574 0 54630 800 6 la_data_in[103]
port 122 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 la_data_in[104]
port 123 nsew signal input
rlabel metal2 s 55402 0 55458 800 6 la_data_in[105]
port 124 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_data_in[106]
port 125 nsew signal input
rlabel metal2 s 56138 0 56194 800 6 la_data_in[107]
port 126 nsew signal input
rlabel metal2 s 56506 0 56562 800 6 la_data_in[108]
port 127 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[109]
port 128 nsew signal input
rlabel metal2 s 17866 0 17922 800 6 la_data_in[10]
port 129 nsew signal input
rlabel metal2 s 57334 0 57390 800 6 la_data_in[110]
port 130 nsew signal input
rlabel metal2 s 57702 0 57758 800 6 la_data_in[111]
port 131 nsew signal input
rlabel metal2 s 58162 0 58218 800 6 la_data_in[112]
port 132 nsew signal input
rlabel metal2 s 58530 0 58586 800 6 la_data_in[113]
port 133 nsew signal input
rlabel metal2 s 58898 0 58954 800 6 la_data_in[114]
port 134 nsew signal input
rlabel metal2 s 59266 0 59322 800 6 la_data_in[115]
port 135 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[116]
port 136 nsew signal input
rlabel metal2 s 60094 0 60150 800 6 la_data_in[117]
port 137 nsew signal input
rlabel metal2 s 60462 0 60518 800 6 la_data_in[118]
port 138 nsew signal input
rlabel metal2 s 60922 0 60978 800 6 la_data_in[119]
port 139 nsew signal input
rlabel metal2 s 18234 0 18290 800 6 la_data_in[11]
port 140 nsew signal input
rlabel metal2 s 61290 0 61346 800 6 la_data_in[120]
port 141 nsew signal input
rlabel metal2 s 61658 0 61714 800 6 la_data_in[121]
port 142 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[122]
port 143 nsew signal input
rlabel metal2 s 62486 0 62542 800 6 la_data_in[123]
port 144 nsew signal input
rlabel metal2 s 62854 0 62910 800 6 la_data_in[124]
port 145 nsew signal input
rlabel metal2 s 63222 0 63278 800 6 la_data_in[125]
port 146 nsew signal input
rlabel metal2 s 63682 0 63738 800 6 la_data_in[126]
port 147 nsew signal input
rlabel metal2 s 64050 0 64106 800 6 la_data_in[127]
port 148 nsew signal input
rlabel metal2 s 18694 0 18750 800 6 la_data_in[12]
port 149 nsew signal input
rlabel metal2 s 19062 0 19118 800 6 la_data_in[13]
port 150 nsew signal input
rlabel metal2 s 19430 0 19486 800 6 la_data_in[14]
port 151 nsew signal input
rlabel metal2 s 19798 0 19854 800 6 la_data_in[15]
port 152 nsew signal input
rlabel metal2 s 20258 0 20314 800 6 la_data_in[16]
port 153 nsew signal input
rlabel metal2 s 20626 0 20682 800 6 la_data_in[17]
port 154 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 la_data_in[18]
port 155 nsew signal input
rlabel metal2 s 21454 0 21510 800 6 la_data_in[19]
port 156 nsew signal input
rlabel metal2 s 14278 0 14334 800 6 la_data_in[1]
port 157 nsew signal input
rlabel metal2 s 21822 0 21878 800 6 la_data_in[20]
port 158 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 la_data_in[21]
port 159 nsew signal input
rlabel metal2 s 22558 0 22614 800 6 la_data_in[22]
port 160 nsew signal input
rlabel metal2 s 23018 0 23074 800 6 la_data_in[23]
port 161 nsew signal input
rlabel metal2 s 23386 0 23442 800 6 la_data_in[24]
port 162 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 la_data_in[25]
port 163 nsew signal input
rlabel metal2 s 24214 0 24270 800 6 la_data_in[26]
port 164 nsew signal input
rlabel metal2 s 24582 0 24638 800 6 la_data_in[27]
port 165 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 la_data_in[28]
port 166 nsew signal input
rlabel metal2 s 25318 0 25374 800 6 la_data_in[29]
port 167 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 la_data_in[2]
port 168 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 la_data_in[30]
port 169 nsew signal input
rlabel metal2 s 26146 0 26202 800 6 la_data_in[31]
port 170 nsew signal input
rlabel metal2 s 26514 0 26570 800 6 la_data_in[32]
port 171 nsew signal input
rlabel metal2 s 26974 0 27030 800 6 la_data_in[33]
port 172 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 la_data_in[34]
port 173 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 la_data_in[35]
port 174 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[36]
port 175 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 la_data_in[37]
port 176 nsew signal input
rlabel metal2 s 28906 0 28962 800 6 la_data_in[38]
port 177 nsew signal input
rlabel metal2 s 29274 0 29330 800 6 la_data_in[39]
port 178 nsew signal input
rlabel metal2 s 15106 0 15162 800 6 la_data_in[3]
port 179 nsew signal input
rlabel metal2 s 29734 0 29790 800 6 la_data_in[40]
port 180 nsew signal input
rlabel metal2 s 30102 0 30158 800 6 la_data_in[41]
port 181 nsew signal input
rlabel metal2 s 30470 0 30526 800 6 la_data_in[42]
port 182 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 la_data_in[43]
port 183 nsew signal input
rlabel metal2 s 31298 0 31354 800 6 la_data_in[44]
port 184 nsew signal input
rlabel metal2 s 31666 0 31722 800 6 la_data_in[45]
port 185 nsew signal input
rlabel metal2 s 32034 0 32090 800 6 la_data_in[46]
port 186 nsew signal input
rlabel metal2 s 32494 0 32550 800 6 la_data_in[47]
port 187 nsew signal input
rlabel metal2 s 32862 0 32918 800 6 la_data_in[48]
port 188 nsew signal input
rlabel metal2 s 33230 0 33286 800 6 la_data_in[49]
port 189 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 la_data_in[4]
port 190 nsew signal input
rlabel metal2 s 33690 0 33746 800 6 la_data_in[50]
port 191 nsew signal input
rlabel metal2 s 34058 0 34114 800 6 la_data_in[51]
port 192 nsew signal input
rlabel metal2 s 34426 0 34482 800 6 la_data_in[52]
port 193 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 la_data_in[53]
port 194 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 la_data_in[54]
port 195 nsew signal input
rlabel metal2 s 35622 0 35678 800 6 la_data_in[55]
port 196 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_data_in[56]
port 197 nsew signal input
rlabel metal2 s 36450 0 36506 800 6 la_data_in[57]
port 198 nsew signal input
rlabel metal2 s 36818 0 36874 800 6 la_data_in[58]
port 199 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_data_in[59]
port 200 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 la_data_in[5]
port 201 nsew signal input
rlabel metal2 s 37554 0 37610 800 6 la_data_in[60]
port 202 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 la_data_in[61]
port 203 nsew signal input
rlabel metal2 s 38382 0 38438 800 6 la_data_in[62]
port 204 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_data_in[63]
port 205 nsew signal input
rlabel metal2 s 39210 0 39266 800 6 la_data_in[64]
port 206 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_data_in[65]
port 207 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[66]
port 208 nsew signal input
rlabel metal2 s 40406 0 40462 800 6 la_data_in[67]
port 209 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[68]
port 210 nsew signal input
rlabel metal2 s 41142 0 41198 800 6 la_data_in[69]
port 211 nsew signal input
rlabel metal2 s 16302 0 16358 800 6 la_data_in[6]
port 212 nsew signal input
rlabel metal2 s 41510 0 41566 800 6 la_data_in[70]
port 213 nsew signal input
rlabel metal2 s 41970 0 42026 800 6 la_data_in[71]
port 214 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_data_in[72]
port 215 nsew signal input
rlabel metal2 s 42706 0 42762 800 6 la_data_in[73]
port 216 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_data_in[74]
port 217 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[75]
port 218 nsew signal input
rlabel metal2 s 43902 0 43958 800 6 la_data_in[76]
port 219 nsew signal input
rlabel metal2 s 44270 0 44326 800 6 la_data_in[77]
port 220 nsew signal input
rlabel metal2 s 44730 0 44786 800 6 la_data_in[78]
port 221 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[79]
port 222 nsew signal input
rlabel metal2 s 16670 0 16726 800 6 la_data_in[7]
port 223 nsew signal input
rlabel metal2 s 45466 0 45522 800 6 la_data_in[80]
port 224 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_data_in[81]
port 225 nsew signal input
rlabel metal2 s 46294 0 46350 800 6 la_data_in[82]
port 226 nsew signal input
rlabel metal2 s 46662 0 46718 800 6 la_data_in[83]
port 227 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 la_data_in[84]
port 228 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 la_data_in[85]
port 229 nsew signal input
rlabel metal2 s 47858 0 47914 800 6 la_data_in[86]
port 230 nsew signal input
rlabel metal2 s 48226 0 48282 800 6 la_data_in[87]
port 231 nsew signal input
rlabel metal2 s 48686 0 48742 800 6 la_data_in[88]
port 232 nsew signal input
rlabel metal2 s 49054 0 49110 800 6 la_data_in[89]
port 233 nsew signal input
rlabel metal2 s 17038 0 17094 800 6 la_data_in[8]
port 234 nsew signal input
rlabel metal2 s 49422 0 49478 800 6 la_data_in[90]
port 235 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[91]
port 236 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 la_data_in[92]
port 237 nsew signal input
rlabel metal2 s 50618 0 50674 800 6 la_data_in[93]
port 238 nsew signal input
rlabel metal2 s 50986 0 51042 800 6 la_data_in[94]
port 239 nsew signal input
rlabel metal2 s 51446 0 51502 800 6 la_data_in[95]
port 240 nsew signal input
rlabel metal2 s 51814 0 51870 800 6 la_data_in[96]
port 241 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_data_in[97]
port 242 nsew signal input
rlabel metal2 s 52642 0 52698 800 6 la_data_in[98]
port 243 nsew signal input
rlabel metal2 s 53010 0 53066 800 6 la_data_in[99]
port 244 nsew signal input
rlabel metal2 s 17498 0 17554 800 6 la_data_in[9]
port 245 nsew signal input
rlabel metal2 s 14094 0 14150 800 6 la_data_out[0]
port 246 nsew signal output
rlabel metal2 s 53562 0 53618 800 6 la_data_out[100]
port 247 nsew signal output
rlabel metal2 s 53930 0 53986 800 6 la_data_out[101]
port 248 nsew signal output
rlabel metal2 s 54298 0 54354 800 6 la_data_out[102]
port 249 nsew signal output
rlabel metal2 s 54666 0 54722 800 6 la_data_out[103]
port 250 nsew signal output
rlabel metal2 s 55126 0 55182 800 6 la_data_out[104]
port 251 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[105]
port 252 nsew signal output
rlabel metal2 s 55862 0 55918 800 6 la_data_out[106]
port 253 nsew signal output
rlabel metal2 s 56322 0 56378 800 6 la_data_out[107]
port 254 nsew signal output
rlabel metal2 s 56690 0 56746 800 6 la_data_out[108]
port 255 nsew signal output
rlabel metal2 s 57058 0 57114 800 6 la_data_out[109]
port 256 nsew signal output
rlabel metal2 s 17958 0 18014 800 6 la_data_out[10]
port 257 nsew signal output
rlabel metal2 s 57426 0 57482 800 6 la_data_out[110]
port 258 nsew signal output
rlabel metal2 s 57886 0 57942 800 6 la_data_out[111]
port 259 nsew signal output
rlabel metal2 s 58254 0 58310 800 6 la_data_out[112]
port 260 nsew signal output
rlabel metal2 s 58622 0 58678 800 6 la_data_out[113]
port 261 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[114]
port 262 nsew signal output
rlabel metal2 s 59450 0 59506 800 6 la_data_out[115]
port 263 nsew signal output
rlabel metal2 s 59818 0 59874 800 6 la_data_out[116]
port 264 nsew signal output
rlabel metal2 s 60186 0 60242 800 6 la_data_out[117]
port 265 nsew signal output
rlabel metal2 s 60646 0 60702 800 6 la_data_out[118]
port 266 nsew signal output
rlabel metal2 s 61014 0 61070 800 6 la_data_out[119]
port 267 nsew signal output
rlabel metal2 s 18418 0 18474 800 6 la_data_out[11]
port 268 nsew signal output
rlabel metal2 s 61382 0 61438 800 6 la_data_out[120]
port 269 nsew signal output
rlabel metal2 s 61842 0 61898 800 6 la_data_out[121]
port 270 nsew signal output
rlabel metal2 s 62210 0 62266 800 6 la_data_out[122]
port 271 nsew signal output
rlabel metal2 s 62578 0 62634 800 6 la_data_out[123]
port 272 nsew signal output
rlabel metal2 s 62946 0 63002 800 6 la_data_out[124]
port 273 nsew signal output
rlabel metal2 s 63406 0 63462 800 6 la_data_out[125]
port 274 nsew signal output
rlabel metal2 s 63774 0 63830 800 6 la_data_out[126]
port 275 nsew signal output
rlabel metal2 s 64142 0 64198 800 6 la_data_out[127]
port 276 nsew signal output
rlabel metal2 s 18786 0 18842 800 6 la_data_out[12]
port 277 nsew signal output
rlabel metal2 s 19154 0 19210 800 6 la_data_out[13]
port 278 nsew signal output
rlabel metal2 s 19614 0 19670 800 6 la_data_out[14]
port 279 nsew signal output
rlabel metal2 s 19982 0 20038 800 6 la_data_out[15]
port 280 nsew signal output
rlabel metal2 s 20350 0 20406 800 6 la_data_out[16]
port 281 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 la_data_out[17]
port 282 nsew signal output
rlabel metal2 s 21178 0 21234 800 6 la_data_out[18]
port 283 nsew signal output
rlabel metal2 s 21546 0 21602 800 6 la_data_out[19]
port 284 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 la_data_out[1]
port 285 nsew signal output
rlabel metal2 s 21914 0 21970 800 6 la_data_out[20]
port 286 nsew signal output
rlabel metal2 s 22374 0 22430 800 6 la_data_out[21]
port 287 nsew signal output
rlabel metal2 s 22742 0 22798 800 6 la_data_out[22]
port 288 nsew signal output
rlabel metal2 s 23110 0 23166 800 6 la_data_out[23]
port 289 nsew signal output
rlabel metal2 s 23478 0 23534 800 6 la_data_out[24]
port 290 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 la_data_out[25]
port 291 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 la_data_out[26]
port 292 nsew signal output
rlabel metal2 s 24674 0 24730 800 6 la_data_out[27]
port 293 nsew signal output
rlabel metal2 s 25134 0 25190 800 6 la_data_out[28]
port 294 nsew signal output
rlabel metal2 s 25502 0 25558 800 6 la_data_out[29]
port 295 nsew signal output
rlabel metal2 s 14830 0 14886 800 6 la_data_out[2]
port 296 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 la_data_out[30]
port 297 nsew signal output
rlabel metal2 s 26330 0 26386 800 6 la_data_out[31]
port 298 nsew signal output
rlabel metal2 s 26698 0 26754 800 6 la_data_out[32]
port 299 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 la_data_out[33]
port 300 nsew signal output
rlabel metal2 s 27434 0 27490 800 6 la_data_out[34]
port 301 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 la_data_out[35]
port 302 nsew signal output
rlabel metal2 s 28262 0 28318 800 6 la_data_out[36]
port 303 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 la_data_out[37]
port 304 nsew signal output
rlabel metal2 s 29090 0 29146 800 6 la_data_out[38]
port 305 nsew signal output
rlabel metal2 s 29458 0 29514 800 6 la_data_out[39]
port 306 nsew signal output
rlabel metal2 s 15198 0 15254 800 6 la_data_out[3]
port 307 nsew signal output
rlabel metal2 s 29826 0 29882 800 6 la_data_out[40]
port 308 nsew signal output
rlabel metal2 s 30194 0 30250 800 6 la_data_out[41]
port 309 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 la_data_out[42]
port 310 nsew signal output
rlabel metal2 s 31022 0 31078 800 6 la_data_out[43]
port 311 nsew signal output
rlabel metal2 s 31390 0 31446 800 6 la_data_out[44]
port 312 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 la_data_out[45]
port 313 nsew signal output
rlabel metal2 s 32218 0 32274 800 6 la_data_out[46]
port 314 nsew signal output
rlabel metal2 s 32586 0 32642 800 6 la_data_out[47]
port 315 nsew signal output
rlabel metal2 s 32954 0 33010 800 6 la_data_out[48]
port 316 nsew signal output
rlabel metal2 s 33414 0 33470 800 6 la_data_out[49]
port 317 nsew signal output
rlabel metal2 s 15658 0 15714 800 6 la_data_out[4]
port 318 nsew signal output
rlabel metal2 s 33782 0 33838 800 6 la_data_out[50]
port 319 nsew signal output
rlabel metal2 s 34150 0 34206 800 6 la_data_out[51]
port 320 nsew signal output
rlabel metal2 s 34610 0 34666 800 6 la_data_out[52]
port 321 nsew signal output
rlabel metal2 s 34978 0 35034 800 6 la_data_out[53]
port 322 nsew signal output
rlabel metal2 s 35346 0 35402 800 6 la_data_out[54]
port 323 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 la_data_out[55]
port 324 nsew signal output
rlabel metal2 s 36174 0 36230 800 6 la_data_out[56]
port 325 nsew signal output
rlabel metal2 s 36542 0 36598 800 6 la_data_out[57]
port 326 nsew signal output
rlabel metal2 s 36910 0 36966 800 6 la_data_out[58]
port 327 nsew signal output
rlabel metal2 s 37370 0 37426 800 6 la_data_out[59]
port 328 nsew signal output
rlabel metal2 s 16026 0 16082 800 6 la_data_out[5]
port 329 nsew signal output
rlabel metal2 s 37738 0 37794 800 6 la_data_out[60]
port 330 nsew signal output
rlabel metal2 s 38106 0 38162 800 6 la_data_out[61]
port 331 nsew signal output
rlabel metal2 s 38474 0 38530 800 6 la_data_out[62]
port 332 nsew signal output
rlabel metal2 s 38934 0 38990 800 6 la_data_out[63]
port 333 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[64]
port 334 nsew signal output
rlabel metal2 s 39670 0 39726 800 6 la_data_out[65]
port 335 nsew signal output
rlabel metal2 s 40130 0 40186 800 6 la_data_out[66]
port 336 nsew signal output
rlabel metal2 s 40498 0 40554 800 6 la_data_out[67]
port 337 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[68]
port 338 nsew signal output
rlabel metal2 s 41326 0 41382 800 6 la_data_out[69]
port 339 nsew signal output
rlabel metal2 s 16394 0 16450 800 6 la_data_out[6]
port 340 nsew signal output
rlabel metal2 s 41694 0 41750 800 6 la_data_out[70]
port 341 nsew signal output
rlabel metal2 s 42062 0 42118 800 6 la_data_out[71]
port 342 nsew signal output
rlabel metal2 s 42430 0 42486 800 6 la_data_out[72]
port 343 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[73]
port 344 nsew signal output
rlabel metal2 s 43258 0 43314 800 6 la_data_out[74]
port 345 nsew signal output
rlabel metal2 s 43626 0 43682 800 6 la_data_out[75]
port 346 nsew signal output
rlabel metal2 s 44086 0 44142 800 6 la_data_out[76]
port 347 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 la_data_out[77]
port 348 nsew signal output
rlabel metal2 s 44822 0 44878 800 6 la_data_out[78]
port 349 nsew signal output
rlabel metal2 s 45190 0 45246 800 6 la_data_out[79]
port 350 nsew signal output
rlabel metal2 s 16854 0 16910 800 6 la_data_out[7]
port 351 nsew signal output
rlabel metal2 s 45650 0 45706 800 6 la_data_out[80]
port 352 nsew signal output
rlabel metal2 s 46018 0 46074 800 6 la_data_out[81]
port 353 nsew signal output
rlabel metal2 s 46386 0 46442 800 6 la_data_out[82]
port 354 nsew signal output
rlabel metal2 s 46846 0 46902 800 6 la_data_out[83]
port 355 nsew signal output
rlabel metal2 s 47214 0 47270 800 6 la_data_out[84]
port 356 nsew signal output
rlabel metal2 s 47582 0 47638 800 6 la_data_out[85]
port 357 nsew signal output
rlabel metal2 s 47950 0 48006 800 6 la_data_out[86]
port 358 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 la_data_out[87]
port 359 nsew signal output
rlabel metal2 s 48778 0 48834 800 6 la_data_out[88]
port 360 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 la_data_out[89]
port 361 nsew signal output
rlabel metal2 s 17222 0 17278 800 6 la_data_out[8]
port 362 nsew signal output
rlabel metal2 s 49606 0 49662 800 6 la_data_out[90]
port 363 nsew signal output
rlabel metal2 s 49974 0 50030 800 6 la_data_out[91]
port 364 nsew signal output
rlabel metal2 s 50342 0 50398 800 6 la_data_out[92]
port 365 nsew signal output
rlabel metal2 s 50710 0 50766 800 6 la_data_out[93]
port 366 nsew signal output
rlabel metal2 s 51170 0 51226 800 6 la_data_out[94]
port 367 nsew signal output
rlabel metal2 s 51538 0 51594 800 6 la_data_out[95]
port 368 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[96]
port 369 nsew signal output
rlabel metal2 s 52366 0 52422 800 6 la_data_out[97]
port 370 nsew signal output
rlabel metal2 s 52734 0 52790 800 6 la_data_out[98]
port 371 nsew signal output
rlabel metal2 s 53102 0 53158 800 6 la_data_out[99]
port 372 nsew signal output
rlabel metal2 s 17590 0 17646 800 6 la_data_out[9]
port 373 nsew signal output
rlabel metal2 s 14186 0 14242 800 6 la_oenb[0]
port 374 nsew signal input
rlabel metal2 s 53654 0 53710 800 6 la_oenb[100]
port 375 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[101]
port 376 nsew signal input
rlabel metal2 s 54482 0 54538 800 6 la_oenb[102]
port 377 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[103]
port 378 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_oenb[104]
port 379 nsew signal input
rlabel metal2 s 55586 0 55642 800 6 la_oenb[105]
port 380 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_oenb[106]
port 381 nsew signal input
rlabel metal2 s 56414 0 56470 800 6 la_oenb[107]
port 382 nsew signal input
rlabel metal2 s 56782 0 56838 800 6 la_oenb[108]
port 383 nsew signal input
rlabel metal2 s 57242 0 57298 800 6 la_oenb[109]
port 384 nsew signal input
rlabel metal2 s 18142 0 18198 800 6 la_oenb[10]
port 385 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[110]
port 386 nsew signal input
rlabel metal2 s 57978 0 58034 800 6 la_oenb[111]
port 387 nsew signal input
rlabel metal2 s 58346 0 58402 800 6 la_oenb[112]
port 388 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_oenb[113]
port 389 nsew signal input
rlabel metal2 s 59174 0 59230 800 6 la_oenb[114]
port 390 nsew signal input
rlabel metal2 s 59542 0 59598 800 6 la_oenb[115]
port 391 nsew signal input
rlabel metal2 s 60002 0 60058 800 6 la_oenb[116]
port 392 nsew signal input
rlabel metal2 s 60370 0 60426 800 6 la_oenb[117]
port 393 nsew signal input
rlabel metal2 s 60738 0 60794 800 6 la_oenb[118]
port 394 nsew signal input
rlabel metal2 s 61106 0 61162 800 6 la_oenb[119]
port 395 nsew signal input
rlabel metal2 s 18510 0 18566 800 6 la_oenb[11]
port 396 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 la_oenb[120]
port 397 nsew signal input
rlabel metal2 s 61934 0 61990 800 6 la_oenb[121]
port 398 nsew signal input
rlabel metal2 s 62302 0 62358 800 6 la_oenb[122]
port 399 nsew signal input
rlabel metal2 s 62762 0 62818 800 6 la_oenb[123]
port 400 nsew signal input
rlabel metal2 s 63130 0 63186 800 6 la_oenb[124]
port 401 nsew signal input
rlabel metal2 s 63498 0 63554 800 6 la_oenb[125]
port 402 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[126]
port 403 nsew signal input
rlabel metal2 s 64326 0 64382 800 6 la_oenb[127]
port 404 nsew signal input
rlabel metal2 s 18878 0 18934 800 6 la_oenb[12]
port 405 nsew signal input
rlabel metal2 s 19338 0 19394 800 6 la_oenb[13]
port 406 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la_oenb[14]
port 407 nsew signal input
rlabel metal2 s 20074 0 20130 800 6 la_oenb[15]
port 408 nsew signal input
rlabel metal2 s 20534 0 20590 800 6 la_oenb[16]
port 409 nsew signal input
rlabel metal2 s 20902 0 20958 800 6 la_oenb[17]
port 410 nsew signal input
rlabel metal2 s 21270 0 21326 800 6 la_oenb[18]
port 411 nsew signal input
rlabel metal2 s 21638 0 21694 800 6 la_oenb[19]
port 412 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 la_oenb[1]
port 413 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 la_oenb[20]
port 414 nsew signal input
rlabel metal2 s 22466 0 22522 800 6 la_oenb[21]
port 415 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 la_oenb[22]
port 416 nsew signal input
rlabel metal2 s 23294 0 23350 800 6 la_oenb[23]
port 417 nsew signal input
rlabel metal2 s 23662 0 23718 800 6 la_oenb[24]
port 418 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 la_oenb[25]
port 419 nsew signal input
rlabel metal2 s 24398 0 24454 800 6 la_oenb[26]
port 420 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 la_oenb[27]
port 421 nsew signal input
rlabel metal2 s 25226 0 25282 800 6 la_oenb[28]
port 422 nsew signal input
rlabel metal2 s 25594 0 25650 800 6 la_oenb[29]
port 423 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 la_oenb[2]
port 424 nsew signal input
rlabel metal2 s 26054 0 26110 800 6 la_oenb[30]
port 425 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 la_oenb[31]
port 426 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 la_oenb[32]
port 427 nsew signal input
rlabel metal2 s 27250 0 27306 800 6 la_oenb[33]
port 428 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 la_oenb[34]
port 429 nsew signal input
rlabel metal2 s 27986 0 28042 800 6 la_oenb[35]
port 430 nsew signal input
rlabel metal2 s 28354 0 28410 800 6 la_oenb[36]
port 431 nsew signal input
rlabel metal2 s 28814 0 28870 800 6 la_oenb[37]
port 432 nsew signal input
rlabel metal2 s 29182 0 29238 800 6 la_oenb[38]
port 433 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 la_oenb[39]
port 434 nsew signal input
rlabel metal2 s 15382 0 15438 800 6 la_oenb[3]
port 435 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 la_oenb[40]
port 436 nsew signal input
rlabel metal2 s 30378 0 30434 800 6 la_oenb[41]
port 437 nsew signal input
rlabel metal2 s 30746 0 30802 800 6 la_oenb[42]
port 438 nsew signal input
rlabel metal2 s 31114 0 31170 800 6 la_oenb[43]
port 439 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 la_oenb[44]
port 440 nsew signal input
rlabel metal2 s 31942 0 31998 800 6 la_oenb[45]
port 441 nsew signal input
rlabel metal2 s 32310 0 32366 800 6 la_oenb[46]
port 442 nsew signal input
rlabel metal2 s 32770 0 32826 800 6 la_oenb[47]
port 443 nsew signal input
rlabel metal2 s 33138 0 33194 800 6 la_oenb[48]
port 444 nsew signal input
rlabel metal2 s 33506 0 33562 800 6 la_oenb[49]
port 445 nsew signal input
rlabel metal2 s 15750 0 15806 800 6 la_oenb[4]
port 446 nsew signal input
rlabel metal2 s 33874 0 33930 800 6 la_oenb[50]
port 447 nsew signal input
rlabel metal2 s 34334 0 34390 800 6 la_oenb[51]
port 448 nsew signal input
rlabel metal2 s 34702 0 34758 800 6 la_oenb[52]
port 449 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[53]
port 450 nsew signal input
rlabel metal2 s 35530 0 35586 800 6 la_oenb[54]
port 451 nsew signal input
rlabel metal2 s 35898 0 35954 800 6 la_oenb[55]
port 452 nsew signal input
rlabel metal2 s 36266 0 36322 800 6 la_oenb[56]
port 453 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_oenb[57]
port 454 nsew signal input
rlabel metal2 s 37094 0 37150 800 6 la_oenb[58]
port 455 nsew signal input
rlabel metal2 s 37462 0 37518 800 6 la_oenb[59]
port 456 nsew signal input
rlabel metal2 s 16118 0 16174 800 6 la_oenb[5]
port 457 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[60]
port 458 nsew signal input
rlabel metal2 s 38290 0 38346 800 6 la_oenb[61]
port 459 nsew signal input
rlabel metal2 s 38658 0 38714 800 6 la_oenb[62]
port 460 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_oenb[63]
port 461 nsew signal input
rlabel metal2 s 39486 0 39542 800 6 la_oenb[64]
port 462 nsew signal input
rlabel metal2 s 39854 0 39910 800 6 la_oenb[65]
port 463 nsew signal input
rlabel metal2 s 40222 0 40278 800 6 la_oenb[66]
port 464 nsew signal input
rlabel metal2 s 40590 0 40646 800 6 la_oenb[67]
port 465 nsew signal input
rlabel metal2 s 41050 0 41106 800 6 la_oenb[68]
port 466 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[69]
port 467 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 la_oenb[6]
port 468 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 la_oenb[70]
port 469 nsew signal input
rlabel metal2 s 42246 0 42302 800 6 la_oenb[71]
port 470 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_oenb[72]
port 471 nsew signal input
rlabel metal2 s 42982 0 43038 800 6 la_oenb[73]
port 472 nsew signal input
rlabel metal2 s 43350 0 43406 800 6 la_oenb[74]
port 473 nsew signal input
rlabel metal2 s 43810 0 43866 800 6 la_oenb[75]
port 474 nsew signal input
rlabel metal2 s 44178 0 44234 800 6 la_oenb[76]
port 475 nsew signal input
rlabel metal2 s 44546 0 44602 800 6 la_oenb[77]
port 476 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[78]
port 477 nsew signal input
rlabel metal2 s 45374 0 45430 800 6 la_oenb[79]
port 478 nsew signal input
rlabel metal2 s 16946 0 17002 800 6 la_oenb[7]
port 479 nsew signal input
rlabel metal2 s 45742 0 45798 800 6 la_oenb[80]
port 480 nsew signal input
rlabel metal2 s 46110 0 46166 800 6 la_oenb[81]
port 481 nsew signal input
rlabel metal2 s 46570 0 46626 800 6 la_oenb[82]
port 482 nsew signal input
rlabel metal2 s 46938 0 46994 800 6 la_oenb[83]
port 483 nsew signal input
rlabel metal2 s 47306 0 47362 800 6 la_oenb[84]
port 484 nsew signal input
rlabel metal2 s 47766 0 47822 800 6 la_oenb[85]
port 485 nsew signal input
rlabel metal2 s 48134 0 48190 800 6 la_oenb[86]
port 486 nsew signal input
rlabel metal2 s 48502 0 48558 800 6 la_oenb[87]
port 487 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_oenb[88]
port 488 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 la_oenb[89]
port 489 nsew signal input
rlabel metal2 s 17314 0 17370 800 6 la_oenb[8]
port 490 nsew signal input
rlabel metal2 s 49698 0 49754 800 6 la_oenb[90]
port 491 nsew signal input
rlabel metal2 s 50066 0 50122 800 6 la_oenb[91]
port 492 nsew signal input
rlabel metal2 s 50526 0 50582 800 6 la_oenb[92]
port 493 nsew signal input
rlabel metal2 s 50894 0 50950 800 6 la_oenb[93]
port 494 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[94]
port 495 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_oenb[95]
port 496 nsew signal input
rlabel metal2 s 52090 0 52146 800 6 la_oenb[96]
port 497 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_oenb[97]
port 498 nsew signal input
rlabel metal2 s 52826 0 52882 800 6 la_oenb[98]
port 499 nsew signal input
rlabel metal2 s 53286 0 53342 800 6 la_oenb[99]
port 500 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 la_oenb[9]
port 501 nsew signal input
rlabel metal4 s 4208 2128 4528 64784 6 vccd1
port 502 nsew power input
rlabel metal4 s 34928 2128 35248 64784 6 vccd1
port 502 nsew power input
rlabel metal4 s 19568 2128 19888 64784 6 vssd1
port 503 nsew ground input
rlabel metal4 s 50288 2128 50608 64784 6 vssd1
port 503 nsew ground input
rlabel metal2 s 18 0 74 800 6 wb_clk_i
port 504 nsew signal input
rlabel metal2 s 110 0 166 800 6 wb_rst_i
port 505 nsew signal input
rlabel metal2 s 202 0 258 800 6 wbs_ack_o
port 506 nsew signal output
rlabel metal2 s 754 0 810 800 6 wbs_adr_i[0]
port 507 nsew signal input
rlabel metal2 s 5262 0 5318 800 6 wbs_adr_i[10]
port 508 nsew signal input
rlabel metal2 s 5630 0 5686 800 6 wbs_adr_i[11]
port 509 nsew signal input
rlabel metal2 s 5998 0 6054 800 6 wbs_adr_i[12]
port 510 nsew signal input
rlabel metal2 s 6458 0 6514 800 6 wbs_adr_i[13]
port 511 nsew signal input
rlabel metal2 s 6826 0 6882 800 6 wbs_adr_i[14]
port 512 nsew signal input
rlabel metal2 s 7194 0 7250 800 6 wbs_adr_i[15]
port 513 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[16]
port 514 nsew signal input
rlabel metal2 s 8022 0 8078 800 6 wbs_adr_i[17]
port 515 nsew signal input
rlabel metal2 s 8390 0 8446 800 6 wbs_adr_i[18]
port 516 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_adr_i[19]
port 517 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_adr_i[1]
port 518 nsew signal input
rlabel metal2 s 9218 0 9274 800 6 wbs_adr_i[20]
port 519 nsew signal input
rlabel metal2 s 9586 0 9642 800 6 wbs_adr_i[21]
port 520 nsew signal input
rlabel metal2 s 9954 0 10010 800 6 wbs_adr_i[22]
port 521 nsew signal input
rlabel metal2 s 10322 0 10378 800 6 wbs_adr_i[23]
port 522 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_adr_i[24]
port 523 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[25]
port 524 nsew signal input
rlabel metal2 s 11518 0 11574 800 6 wbs_adr_i[26]
port 525 nsew signal input
rlabel metal2 s 11978 0 12034 800 6 wbs_adr_i[27]
port 526 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_adr_i[28]
port 527 nsew signal input
rlabel metal2 s 12714 0 12770 800 6 wbs_adr_i[29]
port 528 nsew signal input
rlabel metal2 s 1858 0 1914 800 6 wbs_adr_i[2]
port 529 nsew signal input
rlabel metal2 s 13174 0 13230 800 6 wbs_adr_i[30]
port 530 nsew signal input
rlabel metal2 s 13542 0 13598 800 6 wbs_adr_i[31]
port 531 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_adr_i[3]
port 532 nsew signal input
rlabel metal2 s 2870 0 2926 800 6 wbs_adr_i[4]
port 533 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_adr_i[5]
port 534 nsew signal input
rlabel metal2 s 3698 0 3754 800 6 wbs_adr_i[6]
port 535 nsew signal input
rlabel metal2 s 4066 0 4122 800 6 wbs_adr_i[7]
port 536 nsew signal input
rlabel metal2 s 4434 0 4490 800 6 wbs_adr_i[8]
port 537 nsew signal input
rlabel metal2 s 4802 0 4858 800 6 wbs_adr_i[9]
port 538 nsew signal input
rlabel metal2 s 386 0 442 800 6 wbs_cyc_i
port 539 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_dat_i[0]
port 540 nsew signal input
rlabel metal2 s 5354 0 5410 800 6 wbs_dat_i[10]
port 541 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[11]
port 542 nsew signal input
rlabel metal2 s 6182 0 6238 800 6 wbs_dat_i[12]
port 543 nsew signal input
rlabel metal2 s 6550 0 6606 800 6 wbs_dat_i[13]
port 544 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[14]
port 545 nsew signal input
rlabel metal2 s 7378 0 7434 800 6 wbs_dat_i[15]
port 546 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 wbs_dat_i[16]
port 547 nsew signal input
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_i[17]
port 548 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_dat_i[18]
port 549 nsew signal input
rlabel metal2 s 8942 0 8998 800 6 wbs_dat_i[19]
port 550 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wbs_dat_i[1]
port 551 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_dat_i[20]
port 552 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[21]
port 553 nsew signal input
rlabel metal2 s 10138 0 10194 800 6 wbs_dat_i[22]
port 554 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[23]
port 555 nsew signal input
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_i[24]
port 556 nsew signal input
rlabel metal2 s 11242 0 11298 800 6 wbs_dat_i[25]
port 557 nsew signal input
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_i[26]
port 558 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_dat_i[27]
port 559 nsew signal input
rlabel metal2 s 12438 0 12494 800 6 wbs_dat_i[28]
port 560 nsew signal input
rlabel metal2 s 12898 0 12954 800 6 wbs_dat_i[29]
port 561 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 wbs_dat_i[2]
port 562 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[30]
port 563 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_dat_i[31]
port 564 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_i[3]
port 565 nsew signal input
rlabel metal2 s 2962 0 3018 800 6 wbs_dat_i[4]
port 566 nsew signal input
rlabel metal2 s 3422 0 3478 800 6 wbs_dat_i[5]
port 567 nsew signal input
rlabel metal2 s 3790 0 3846 800 6 wbs_dat_i[6]
port 568 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_dat_i[7]
port 569 nsew signal input
rlabel metal2 s 4618 0 4674 800 6 wbs_dat_i[8]
port 570 nsew signal input
rlabel metal2 s 4986 0 5042 800 6 wbs_dat_i[9]
port 571 nsew signal input
rlabel metal2 s 1030 0 1086 800 6 wbs_dat_o[0]
port 572 nsew signal output
rlabel metal2 s 5538 0 5594 800 6 wbs_dat_o[10]
port 573 nsew signal output
rlabel metal2 s 5906 0 5962 800 6 wbs_dat_o[11]
port 574 nsew signal output
rlabel metal2 s 6274 0 6330 800 6 wbs_dat_o[12]
port 575 nsew signal output
rlabel metal2 s 6642 0 6698 800 6 wbs_dat_o[13]
port 576 nsew signal output
rlabel metal2 s 7102 0 7158 800 6 wbs_dat_o[14]
port 577 nsew signal output
rlabel metal2 s 7470 0 7526 800 6 wbs_dat_o[15]
port 578 nsew signal output
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_o[16]
port 579 nsew signal output
rlabel metal2 s 8298 0 8354 800 6 wbs_dat_o[17]
port 580 nsew signal output
rlabel metal2 s 8666 0 8722 800 6 wbs_dat_o[18]
port 581 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[19]
port 582 nsew signal output
rlabel metal2 s 1582 0 1638 800 6 wbs_dat_o[1]
port 583 nsew signal output
rlabel metal2 s 9402 0 9458 800 6 wbs_dat_o[20]
port 584 nsew signal output
rlabel metal2 s 9862 0 9918 800 6 wbs_dat_o[21]
port 585 nsew signal output
rlabel metal2 s 10230 0 10286 800 6 wbs_dat_o[22]
port 586 nsew signal output
rlabel metal2 s 10598 0 10654 800 6 wbs_dat_o[23]
port 587 nsew signal output
rlabel metal2 s 11058 0 11114 800 6 wbs_dat_o[24]
port 588 nsew signal output
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_o[25]
port 589 nsew signal output
rlabel metal2 s 11794 0 11850 800 6 wbs_dat_o[26]
port 590 nsew signal output
rlabel metal2 s 12162 0 12218 800 6 wbs_dat_o[27]
port 591 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[28]
port 592 nsew signal output
rlabel metal2 s 12990 0 13046 800 6 wbs_dat_o[29]
port 593 nsew signal output
rlabel metal2 s 2042 0 2098 800 6 wbs_dat_o[2]
port 594 nsew signal output
rlabel metal2 s 13358 0 13414 800 6 wbs_dat_o[30]
port 595 nsew signal output
rlabel metal2 s 13818 0 13874 800 6 wbs_dat_o[31]
port 596 nsew signal output
rlabel metal2 s 2594 0 2650 800 6 wbs_dat_o[3]
port 597 nsew signal output
rlabel metal2 s 3146 0 3202 800 6 wbs_dat_o[4]
port 598 nsew signal output
rlabel metal2 s 3514 0 3570 800 6 wbs_dat_o[5]
port 599 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 wbs_dat_o[6]
port 600 nsew signal output
rlabel metal2 s 4342 0 4398 800 6 wbs_dat_o[7]
port 601 nsew signal output
rlabel metal2 s 4710 0 4766 800 6 wbs_dat_o[8]
port 602 nsew signal output
rlabel metal2 s 5078 0 5134 800 6 wbs_dat_o[9]
port 603 nsew signal output
rlabel metal2 s 1122 0 1178 800 6 wbs_sel_i[0]
port 604 nsew signal input
rlabel metal2 s 1674 0 1730 800 6 wbs_sel_i[1]
port 605 nsew signal input
rlabel metal2 s 2226 0 2282 800 6 wbs_sel_i[2]
port 606 nsew signal input
rlabel metal2 s 2778 0 2834 800 6 wbs_sel_i[3]
port 607 nsew signal input
rlabel metal2 s 478 0 534 800 6 wbs_stb_i
port 608 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_we_i
port 609 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 64841 66985
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9189310
string GDS_FILE /home/proppy/src/caravel_tutorial/caravel_user_project/openlane/user_proj_example/runs/user_proj_example/results/finishing/user_proj_example.magic.gds
string GDS_START 1003898
<< end >>

